`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: BU
// Engineer: Josh Wildey
// 
// Create Date:    14:36:25 03/17/2018 
// Module Name:    i2c_master 
// Project Name:   PiCamera
// Target Devices: Nexys3 Spartan 6
// Revision 0.01 - File Created
// Description: 
//
// This module will act as a I2C Master Controller
//
//////////////////////////////////////////////////////////////////////////////////
module i2c_master(
	input wire clk,
	input wire rst
    );


endmodule
