`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: BU
// Engineer: Josh Wildey
// 
// Create Date:    14:31:26 04/07/2018 
// Module Name:    keyboard_controller 
// Project Name: Lab 2 - Peripheral and Processor Integration with I/O
// Target Devices: Nexys3 Spartan 6
// Revision 0.01 - File Created
//
//////////////////////////////////////////////////////////////////////////////////
module keyboard_controller(
	input wire       clk,  // Clock from keyboard
	input wire       data, // Data from keyboard
	output reg [7:0] key   // Key pressed on keyboard
   );


endmodule
