`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: J. Wildey
// Module Name: Question 4 a
// Description: Structural verilog
//////////////////////////////////////////////////////////////////////////////////
module question4a(
    input  [3:0] in,
    output [2:0] out
    );


endmodule
